module alu()

endmodule